* Extracted by KLayout

.SUBCKT TOP Q A VSS
M$1 Q A VSS VSS NCHOR1EX L=1U W=2U AS=4P AD=4P PS=8U PD=8U
M$2 Q A \$5 \$5 PCHOR1EX L=1U W=2U AS=4P AD=4P PS=8U PD=8U
.ENDS TOP
